module basic_string;
  string name = "DHANASAKAR";
  
  initial begin
    $display("string name is %s",name.tolower());
  end
endmodule 
