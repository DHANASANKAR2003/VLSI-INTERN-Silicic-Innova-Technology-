module basic_string;
  string name = "DHANASANKAR";
  
  initial begin
    $display("string name is %s",name);
  end
endmodule 
