module basic_string;
  string name = "dhanasankar";
  
  initial begin
    $display("string name is %s",name.toupper());
  end
endmodule 
