`ifndef HA_INTERFACE_SV
`define HA_INTERFACE_SV
interface ha_interface;
  logic a;
  logic b;
  logic s;
  logic c;
  
  event drv_done;
endinterface

`endif
