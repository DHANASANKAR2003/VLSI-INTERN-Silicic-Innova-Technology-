module top_module(
    output zero
);// Module body starts after semicolon
    assign = 1'b0;

endmodule
