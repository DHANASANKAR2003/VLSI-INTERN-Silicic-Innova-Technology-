module basic_string;
  string name = "DHANASANKAR";
  
  initial begin
    $display("string name is %0d",name.len());
  end
endmodule 
